/* Testbench top with nested program to keep Module separated */


// Top module
module tb_top();
endmodule