/* Register file main including parameter and defines */


// Classes tests
program test_p();
endprogram

class testclass;
    string ln;
    rand tsttype test_sel;
    function new(string name);
        ln = name;
    endfunction
endclass

// Macros if needed